module substractor_module
(
    input logic [3:0] coffee_type,
    input logic total_coins,
    input logic cancel_button,
    output logic change,
    output logic enable_timer
);


endmodule
