module coffee_machine
(
);

endmodule 